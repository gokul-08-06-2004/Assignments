// 10.Part Select Operation
// Extract lower nibble from reg [7:0] bus using bus[3:0].

module question_10;
  
  reg [7:0]bus;
  reg [3:0]lower_nibble;
  
  initial begin
    
    bus=8'b10000010;
    
    lower_nibble=bus[3:0];
    
    $display("%b",bus);
    
    $display("%b",lower_nibble);
    
  end
endmodule
